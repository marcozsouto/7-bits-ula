library verilog;
use verilog.vl_types.all;
entity Full_Subtractor_vlg_vec_tst is
end Full_Subtractor_vlg_vec_tst;
