library verilog;
use verilog.vl_types.all;
entity Seven_Segment_Display_vlg_vec_tst is
end Seven_Segment_Display_vlg_vec_tst;
