library verilog;
use verilog.vl_types.all;
entity And_Mux_vlg_vec_tst is
end And_Mux_vlg_vec_tst;
