library verilog;
use verilog.vl_types.all;
entity ULA_Seven_Segments_output_vlg_vec_tst is
end ULA_Seven_Segments_output_vlg_vec_tst;
