library verilog;
use verilog.vl_types.all;
entity BCD_Conversor_vlg_vec_tst is
end BCD_Conversor_vlg_vec_tst;
