library verilog;
use verilog.vl_types.all;
entity Twos_Complement_vlg_vec_tst is
end Twos_Complement_vlg_vec_tst;
