library verilog;
use verilog.vl_types.all;
entity Subtraction_Overflow_vlg_vec_tst is
end Subtraction_Overflow_vlg_vec_tst;
