library verilog;
use verilog.vl_types.all;
entity Seven_bit_Biggest_Comparator_vlg_vec_tst is
end Seven_bit_Biggest_Comparator_vlg_vec_tst;
