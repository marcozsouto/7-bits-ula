library verilog;
use verilog.vl_types.all;
entity Coversor_Seven_Segments_vlg_vec_tst is
end Coversor_Seven_Segments_vlg_vec_tst;
